
module INT 
#(	parameter Win=XX,					// Input
	parameter Wg= XX	) 					// Crecimiento del dato
  (input signed [XX-1:0] data_in, 	// Input data
   input clk,
   input rst,
   input val_in,  					// Validation input
   output reg val_out,					// Validation output
   output reg signed [XX-1:0] data_out);// Output data
	
	
   always@(posedge clk)

	end
		  
		    
	 
endmodule 