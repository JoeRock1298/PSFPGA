module CIC_pc
#(parameter Win=16, // Input length
  parameter Wg=XX)  // Guard bits

  (input signed [Win-1:0] i_data,  		// Data input
   input clk,
   input rst,
   input val_in,  						// Validation input
   output val_out,						// Validation output
   output signed [Win+Wg-1:0] o_data);	// Data output

	

	
	
	//// Insertar la descripción del modulo
	
	
	endmodule 




