module COMB 
#(parameter Win=XX) // Input length
  (input signed [Win-1:0] data_in,
   input clk,
   input rst,
   input val_in,  					// Validation input
   output reg val_out,					// Validation output
   output reg signed  [XX-1:0] data_out);
	
	//// Insertar la descripción del modulo
	

	
	 
endmodule 
