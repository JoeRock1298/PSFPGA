module RD_CONTROL
(
	input txbusy,
	input start_rd,
	input rst, 
	input clk,
	output txena,
	output load_txregs,
	output shift_txregs,
	output done_rd,
	output [2:0] rd_leds
	);


endmodule 