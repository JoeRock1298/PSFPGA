module R_INT
#(parameter Win=XX)
  (input signed [Win-1:0] data_in,
   input clk,
   input rst,
   input val_in,  					// Validation input
   output reg val_out,					// Validation output
   output reg signed [Win-1:0] data_out);



endmodule
			

   