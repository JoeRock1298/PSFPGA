module WR_CONTROL
(
	input rxrdy,
	input start_wr,
	input rst, 
	input clk,
	output shift_rxregs,
	output load_confregs,
	output done_wr,
	output [2:0] wr_leds
	);


	
endmodule 